module tester(
    x,y,eq
);

input wire eq;
output reg x,y;

initial begin
    x=1;
    y=1;
end

endmodule