module tester(
    x,y,eq
);

input wire eq;
output reg x,y;

initial begin
    x=11;
    y=10;
end

endmodule