module tester(
    A_valor, B_valor, N, n_valor
);

input wire N;
output reg A_valor,B_valor,n_valor;

initial begin
    A_valor=1;
    B_valor=1;
    n_valor=0;
    end
endmodule
