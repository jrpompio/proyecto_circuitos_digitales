module Final_ID(
    m, n, A, B, Z;
);
