module Inicial_ID(
    A, B, M, N
);
in